`ifndef _img1_vh_
`define _img1_vh_
    defparam rom1.INIT_RAM_00 = 256'h000000000000000000000000000000003C3834302C2824201C1814100C080400;
    defparam rom1.INIT_RAM_01 = 256'h1010101010101010101010101010101011111111111011110D04000000000000;
    defparam rom1.INIT_RAM_02 = 256'h0000000000000000040F11111111111111111110101010111111111111111212;
    defparam rom1.INIT_RAM_03 = 256'h101010101010101010101010101010101111111111100E040000000000000000;
    defparam rom1.INIT_RAM_04 = 256'h000000000000000000020F111111111111111111111111111111111111111212;
    defparam rom1.INIT_RAM_05 = 256'h1010101010101010101010111111101011111111100E02000000000000000000;
    defparam rom1.INIT_RAM_06 = 256'h0D0D0D1F1F1F17070000020E1010111111111111111111111111111111111212;
    defparam rom1.INIT_RAM_07 = 256'h10101010101010101111111111111111111111100E02000007070D0D0D141414;
    defparam rom1.INIT_RAM_08 = 256'h0D0D0D1F1F1F1F1F170300020E10111111111111111111111111111111111212;
    defparam rom1.INIT_RAM_09 = 256'h101010101010101011111111111111111110100E0200000607070D0D0D141414;
    defparam rom1.INIT_RAM_0A = 256'h0D0F1D1F1F1F1F1F1F1B0300020E111111111111111111111111111111111112;
    defparam rom1.INIT_RAM_0B = 256'h1010101010101010111111111111111111100E0200000607080C0D0D0D14130E;
    defparam rom1.INIT_RAM_0C = 256'h0D1A1F1F1F1F1F1F1F1F1B0300020F1111111111111111111111111111111111;
    defparam rom1.INIT_RAM_0D = 256'h111010101010101008000000020F1111110E0200000507070B0D0D1214100D0D;
    defparam rom1.INIT_RAM_0E = 256'h111F1F1F1F1F1F1F1F1F1F1F0000021111111110101111111111111111111111;
    defparam rom1.INIT_RAM_0F = 256'h11111010101010100000000000020F110F020000010707090D0D0F14140D0D0D;
    defparam rom1.INIT_RAM_10 = 256'h1A1F1F1F1F1F1F1F1F1F1B030000001111111111111111111111111111111111;
    defparam rom1.INIT_RAM_11 = 256'h11101010101010100000000000000211020000000507070B0D0D1214140D0D0D;
    defparam rom1.INIT_RAM_12 = 256'h1F1F1F1F1F1F1F1F1F1B03000000001111111111111111111111111111111112;
    defparam rom1.INIT_RAM_13 = 256'h10111011101010100000000A11020000000000000507070D0D0D1414140D0D0D;
    defparam rom1.INIT_RAM_14 = 256'h1F1F1F1F1F1F1F1F1F0000000000001111111111111111111111111111111212;
    defparam rom1.INIT_RAM_15 = 256'h10101111111010100200001114110000000000000107070D0D0D1414140D0D0D;
    defparam rom1.INIT_RAM_16 = 256'h1F1F1F1F1F1F1F1F1F1B03000000001111111111111111111111111111111212;
    defparam rom1.INIT_RAM_17 = 256'h10101111111010100E02000211141102000000000005070A0D0D1414140D0D0D;
    defparam rom1.INIT_RAM_18 = 256'h1A1F1F1F1F1F1F1F1F1F1B030000001111111111111111111111111111111111;
    defparam rom1.INIT_RAM_19 = 256'h1010101010101010100C0000000A1411020000000000060707071414140D0D0D;
    defparam rom1.INIT_RAM_1A = 256'h111F1F1F1F1F1F1F1F1F1F1F0000001111111111111111111111111111111111;
    defparam rom1.INIT_RAM_1B = 256'h10101010101010101010040000001414110500000000000607071414140D0D0D;
    defparam rom1.INIT_RAM_1C = 256'h0D1A1F1F1F1F1F1F1F1F1F1F0000001111111111111111111111111111111111;
    defparam rom1.INIT_RAM_1D = 256'h101010101010101010100C000000141413120C040000000007071414130E0E0D;
    defparam rom1.INIT_RAM_1E = 256'h0D0F1D1F1F1F1F1F1F1D10100400000D11111111111111111111111111111111;
    defparam rom1.INIT_RAM_1F = 256'h11111111101010101010100000001414131110100C0400000000141413100F0F;
    defparam rom1.INIT_RAM_20 = 256'h0E0D0F1A1F1F1F1F1B1210100C00000411111111111111111111111111111111;
    defparam rom1.INIT_RAM_21 = 256'h111111111110101010101000000014141311101010100C02000214141311100F;
    defparam rom1.INIT_RAM_22 = 256'h0F0E0E0F131B1B1310100F11120500000D111111111111111111111111111111;
    defparam rom1.INIT_RAM_23 = 256'h11111111101010101010080000001313121211111111100E0209131413121110;
    defparam rom1.INIT_RAM_24 = 256'h100F0F0F10101010100F0E0E1311020004111111111111111111111111111111;
    defparam rom1.INIT_RAM_25 = 256'h10101010100800000000000000000D1112121313131312101011131414131312;
    defparam rom1.INIT_RAM_26 = 256'h11101010101010100F0E0D0D14141400000D1111111111111111111111111111;
    defparam rom1.INIT_RAM_27 = 256'h1010101010000000000000000000041011131414141413111011131414141413;
    defparam rom1.INIT_RAM_28 = 256'h1211111111111111100E0D0D1414140000041111111111111111111111111111;
    defparam rom1.INIT_RAM_29 = 256'h1010111111000000000000000000000C10121313141413121112131414141413;
    defparam rom1.INIT_RAM_2A = 256'h1313131313131313130707070707070000041111111111111111111111111111;
    defparam rom1.INIT_RAM_2B = 256'h1010111111000000080E0200000000020E101112131414131313141414141414;
    defparam rom1.INIT_RAM_2C = 256'h14141414141414141407070707070700000C1111111111111111111111111111;
    defparam rom1.INIT_RAM_2D = 256'h10101111110200000E100E0400000000020E1011131414141414141414141414;
    defparam rom1.INIT_RAM_2E = 256'h1414141414141414140D07070707030004111111111111111111111111111111;
    defparam rom1.INIT_RAM_2F = 256'h10111111110F0200020E0F0F0903000000020E10121313141414141414141414;
    defparam rom1.INIT_RAM_30 = 256'h141414141414141414141414000000020F111111111111111111111111111111;
    defparam rom1.INIT_RAM_31 = 256'h1110111010110E020000070E0D0D07070300020E101112131414141414141414;
    defparam rom1.INIT_RAM_32 = 256'h1414141414141414141414140000020F11111111111111111111111111111111;
    defparam rom1.INIT_RAM_33 = 256'h111110101010100E0200000B0D0D070707000002101011131414141414141414;
    defparam rom1.INIT_RAM_34 = 256'h14141414141414141414140A00020F1111111111111111111111121212121111;
    defparam rom1.INIT_RAM_35 = 256'h11101010101010100E0200010D0D070703000000101011131414141414141414;
    defparam rom1.INIT_RAM_36 = 256'h000000000000000000000000000D111111111111111111111212121212121211;
    defparam rom1.INIT_RAM_37 = 256'h1011101110101010110F020000000000000000000C10111314140A0000000000;
    defparam rom1.INIT_RAM_38 = 256'h0000000000000000000000000411111111111111111111111212121212121211;
    defparam rom1.INIT_RAM_39 = 256'h101011111110101011110F040000000000000000041011131414000000000000;
    defparam rom1.INIT_RAM_3A = 256'h0000000000000000000000000D11111111111111111111111212121212121211;
    defparam rom1.INIT_RAM_3B = 256'h1011111111101010111111110C04000000000000000C101213140A0000000000;
    defparam rom1.INIT_RAM_3C = 256'h14141414141414140A0000001111111111111111111111111212121212121111;
    defparam rom1.INIT_RAM_3D = 256'h111111111110101010101010101011111111110800020E101112141414141414;
    defparam rom1.INIT_RAM_3E = 256'h1414141414141414140000021010101111111111111111111111111111111111;
    defparam rom1.INIT_RAM_3F = 256'h11111111111010101010101010101111111111110000020C1011131414141414;
`endif // _img1_vh_
